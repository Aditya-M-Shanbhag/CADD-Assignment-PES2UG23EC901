module test;
reg[3:0] a;
wire p,d;
od I1 (a,p,d);
initial
begin
a[3] = 1'b0; a[2] = 1'b0; a[1] = 1'b0; a[0] = 1'b0;
#10 a[3] = 1'b0; a[2] = 1'b0; a[1] = 1'b0; a[0] = 1'b1;
#10 a[3] = 1'b0; a[2] = 1'b0; a[1] = 1'b1; a[0] = 1'b0;
#10 a[3] = 1'b0; a[2] = 1'b0; a[1] = 1'b1; a[0] = 1'b1;
#10 a[3] = 1'b0; a[2] = 1'b1; a[1] = 1'b0; a[0] = 1'b0;
#10 a[3] = 1'b0; a[2] = 1'b1; a[1] = 1'b0; a[0] = 1'b1;
#10 a[3] = 1'b0; a[2] = 1'b1; a[1] = 1'b1; a[0] = 1'b0;
#10 a[3] = 1'b0; a[2] = 1'b1; a[1] = 1'b1; a[0] = 1'b1;
#10 a[3] = 1'b1; a[2] = 1'b0; a[1] = 1'b0; a[0] = 1'b0;
#10 a[3] = 1'b1; a[2] = 1'b0; a[1] = 1'b0; a[0] = 1'b1;
#10 a[3] = 1'b1; a[2] = 1'b0; a[1] = 1'b1; a[0] = 1'b0;
#10 a[3] = 1'b1; a[2] = 1'b0; a[1] = 1'b1; a[0] = 1'b1;
#10 a[3] = 1'b1; a[2] = 1'b1; a[1] = 1'b0; a[0] = 1'b0;
#10 a[3] = 1'b1; a[2] = 1'b1; a[1] = 1'b0; a[0] = 1'b1;
#10 a[3] = 1'b1; a[2] = 1'b1; a[1] = 1'b1; a[0] = 1'b0;
#10 a[3] = 1'b1; a[2] = 1'b1; a[1] = 1'b1; a[0] = 1'b1;
end
endmodule
